pipe_test.cir
; test for piping to python
; d_process circuit connections:
; in:
;    zero or more inputs (vector) 
;    clock (single input) the event driver
;    reset (single line)
; out:
;   one or more outputs (vector)
;
; d_process pipe data
;  header (all byte values):
;    version (ox1 for this test)
;    number of input bits (bits from ngspice to external program)
;    number of output bits (bits back to ngspice)
; note: the header must be returned to ngspice as handshake
;  data packets to program:
;    double float: running time of ng spice (unit probably seconds)
;         note time will be negative after a reset.
;    input bits packed in bytes (1 byte for 1 to 8 bits, 2 bytes for 9 to 15..)
;  data returned to ngspice
;    output bits packed in bytes (minimal 1 byte)
; 
; arguments from d_process seem to be passed in lower case while python argv is case sensitive!

*** analysis type ***
.tran 10ns 30us
v1 1 0 DC 1.0
v2 2 0 DC 0.0
v3 3 0 DC -1.0

.model d_osc1 d_osc (cntl_array=[-1.0 0.0 1.0 2.0] 
+                    freq_array=[0.1e6 0.5e6 8.0e6 12.0e6]
+                    rise_delay=40.0e-9 fall_delay=40.0e-9)

a1 1 clk1 d_osc1 
a2 2 enable d_osc1 
a3 3 up_down d_osc1

; test with python, different log files for tracebility
ap0_4 [enable up_down] clk1 null [q1 q2 q3 q4] proc0
.model proc0 d_process (process_file="pytest" process_params=["-v", "--log_file", "first.log", "counter"])

ap1_4 [up_down enable] clk1 null [o1 o2 o3 o4] proc1
.model proc1 d_process (process_file="pytest", process_params=["shifter","-v", "--log_file", "shifter.log]))

ap4_1 [o1] clk1 null [delay_o2] proc2
.model proc2 d_process (process_file="pytest" process_params=["delay", "-vvv", "--log_file", "delay.log"])

; ap4_1a [q1 q2 q3 q4] clk1 null [qzeros] proc3
; .model proc3 d_process (process_file="prog4in1out")

.control
run
edisplay
eprvcd clk1 enable up_down q1 q2 q3 q4 o1 o2 o3 o4 delay_o2 > pipe_test.vcd
shell gtkwave pipe_test.vcd --script nggtk.tcl &
quit
.endc
.end

